



module AES256_enc(

                );




endmodule