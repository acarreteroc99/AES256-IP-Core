

/****** mul.sv ******/

module mul(/*nombre senyales*/);
